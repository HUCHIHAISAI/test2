module mx1
endmodule
