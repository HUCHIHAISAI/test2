module mx1
  input a,b;
  output y;
endmodule
